library ieee;
    use ieee.numeric_std.all;
    use ieee.std_logic_1164.all;

library work;
    use work.easysim_axi_common_pkg.AXI_RESP_OKAY_SLV;


package easysim_axi_pkg is

end package easysim_axi_pkg;


package body easysim_axi_pkg is

end package body easysim_axi_pkg;
